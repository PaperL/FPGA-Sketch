//
// Copyright (c) 2015 University of Cambridge
// All rights reserved.
//
//
//  File:
//        output_port_lookup_cpu_regs.v
//
//  Module:
//        output_port_lookup_cpu_regs
//
//  Description:
//        This file is automatically generated with the registers towards the CPU/Software
//
// This software was developed by
// Stanford University and the University of Cambridge Computer Laboratory
// under National Science Foundation under Grant No. CNS-0855268,
// the University of Cambridge Computer Laboratory under EPSRC INTERNET Project EP/H040536/1 and
// by the University of Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-11-C-0249 ("MRC2"),
// as part of the DARPA MRC research programme.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//

`include "output_port_lookup_cpu_regs_defines.v"
module output_port_lookup_cpu_regs #(
    parameter bit     [31:0] C_BASE_ADDRESS     = 32'h00000000,
    parameter integer        C_S_AXI_DATA_WIDTH = 32,
    parameter integer        C_S_AXI_ADDR_WIDTH = 32
) (
    // General ports
    input      clk,
    input      resetn,
    // Global Registers
    input      cpu_resetn_soft,
    output reg resetn_soft,
    output reg resetn_sync,

    // Register ports
    input      [         `REG_ID_BITS] id_reg,
    input      [    `REG_VERSION_BITS] version_reg,
    output reg [      `REG_RESET_BITS] reset_reg,
    input      [       `REG_FLIP_BITS] ip2cpu_flip_reg,
    output reg [       `REG_FLIP_BITS] cpu2ip_flip_reg,
    input      [      `REG_DEBUG_BITS] ip2cpu_debug_reg,
    output reg [      `REG_DEBUG_BITS] cpu2ip_debug_reg,
    input      [      `REG_PKTIN_BITS] pktin_reg,
    output reg                         pktin_reg_clear,
    input      [     `REG_PKTOUT_BITS] pktout_reg,
    output reg                         pktout_reg_clear,
    input      [    `REG_ICMPOUT_BITS] icmpout_reg,
    output reg                         icmpout_reg_clear,
    input      [  `REG_TGTIPADDR_BITS] ip2cpu_tgtipaddr_reg,
    output reg [  `REG_TGTIPADDR_BITS] cpu2ip_tgtipaddr_reg,
    input      [   `REG_TGTIPOUT_BITS] tgtipout_reg,
    output reg                         tgtipout_reg_clear,
    input      [`REG_TGTIPOUTLST_BITS] tgtipoutlst_reg,
    input      [ `REG_TGTUDPPORT_BITS] ip2cpu_tgtudpport_reg,
    output reg [ `REG_TGTUDPPORT_BITS] cpu2ip_tgtudpport_reg,
    input      [  `REG_TGTUDPCNT_BITS] tgtudpcnt_reg,

    // AXI Lite ports
    input                               S_AXI_ACLK,
    input                               S_AXI_ARESETN,
    input  [  C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
    input                               S_AXI_AWVALID,
    input  [  C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
    input  [C_S_AXI_DATA_WIDTH/8-1 : 0] S_AXI_WSTRB,
    input                               S_AXI_WVALID,
    input                               S_AXI_BREADY,
    input  [  C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
    input                               S_AXI_ARVALID,
    input                               S_AXI_RREADY,
    output                              S_AXI_ARREADY,
    output [  C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
    output [                     1 : 0] S_AXI_RRESP,
    output                              S_AXI_RVALID,
    output                              S_AXI_WREADY,
    output [                     1 : 0] S_AXI_BRESP,
    output                              S_AXI_BVALID,
    output                              S_AXI_AWREADY

);

  // AXI4LITE signals
  reg     [C_S_AXI_ADDR_WIDTH-1 : 0] axi_awaddr;
  reg                                axi_awready;
  reg                                axi_wready;
  reg     [                   1 : 0] axi_bresp;
  reg                                axi_bvalid;
  reg     [C_S_AXI_ADDR_WIDTH-1 : 0] axi_araddr;
  reg                                axi_arready;
  reg     [C_S_AXI_DATA_WIDTH-1 : 0] axi_rdata;
  reg     [                   1 : 0] axi_rresp;
  reg                                axi_rvalid;

  reg                                resetn_sync_d;
  wire                               reg_rden;
  wire                               reg_wren;
  reg     [  C_S_AXI_DATA_WIDTH-1:0] reg_data_out;
  integer                            byte_index;
  reg                                pktin_reg_clear_d;
  reg                                pktout_reg_clear_d;
  reg                                icmpout_reg_clear_d;
  reg                                tgtipout_reg_clear_d;

  // I/O Connections assignments
  assign S_AXI_AWREADY = axi_awready;
  assign S_AXI_WREADY  = axi_wready;
  assign S_AXI_BRESP   = axi_bresp;
  assign S_AXI_BVALID  = axi_bvalid;
  assign S_AXI_ARREADY = axi_arready;
  assign S_AXI_RDATA   = axi_rdata;
  assign S_AXI_RRESP   = axi_rresp;
  assign S_AXI_RVALID  = axi_rvalid;

  //Sample reset (not mandatory, but good practice)
  always @(posedge clk) begin
    if (~resetn) begin
      resetn_sync_d <= 1'b0;
      resetn_sync   <= 1'b0;
    end else begin
      resetn_sync_d <= resetn;
      resetn_sync   <= resetn_sync_d;
    end
  end


  /////////////////////////////////
  ////    PROCESS AXI
  /////////////////////////////////


  //global registers, sampling
  always @(posedge clk) resetn_soft <= #1 cpu_resetn_soft;

  // Implement axi_awready generation
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_awready <= 1'b0;
    end else begin
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID) begin
        // slave is ready to accept write address when
        // there is a valid write address and write data
        // on the write address and data bus. This design
        // expects no outstanding transactions.
        axi_awready <= 1'b1;
      end else begin
        axi_awready <= 1'b0;
      end
    end
  end

  // Implement axi_awaddr latching
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_awaddr <= 0;
    end else begin
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID) begin
        // Write Address latching
        axi_awaddr <= S_AXI_AWADDR ^ C_BASE_ADDRESS;
      end
    end
  end

  // Implement axi_wready generation
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_wready <= 1'b0;
    end else begin
      if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID) begin
        // slave is ready to accept write data when
        // there is a valid write address and write data
        // on the write address and data bus. This design
        // expects no outstanding transactions.
        axi_wready <= 1'b1;
      end else begin
        axi_wready <= 1'b0;
      end
    end
  end

  // Implement write response logic generation
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_bvalid <= 0;
      axi_bresp  <= 2'b0;
    end else begin
      if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID) begin
        // indicates a valid write response is available
        axi_bvalid <= 1'b1;
        axi_bresp  <= 2'b0;  // OKAY response
      end                   // work error responses in future
          else
            begin
        if (S_AXI_BREADY && axi_bvalid)
                //check if bready is asserted while bvalid is high)
                //(there is a possibility that bready is always asserted high)
                begin
          axi_bvalid <= 1'b0;
        end
      end
    end
  end

  // Implement axi_arready generation
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_arready <= 1'b0;
      axi_araddr  <= 32'b0;
    end else begin
      if (~axi_arready && S_AXI_ARVALID) begin
        // indicates that the slave has acceped the valid read address
        // Read address latching
        axi_arready <= 1'b1;
        axi_araddr  <= S_AXI_ARADDR ^ C_BASE_ADDRESS;
      end else begin
        axi_arready <= 1'b0;
      end
    end
  end

  // Implement axi_rvalid generation
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_rvalid <= 0;
      axi_rresp  <= 0;
    end else begin
      if (axi_arready && S_AXI_ARVALID && ~axi_rvalid) begin
        // Valid read data is available at the read data bus
        axi_rvalid <= 1'b1;
        axi_rresp  <= 2'b0;  // OKAY response
      end else if (axi_rvalid && S_AXI_RREADY) begin
        // Read data is accepted by the master
        axi_rvalid <= 1'b0;
      end
    end
  end

  // Implement memory mapped register select and write logic generation
  assign reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;


  /////////////////////////////////
  ////    WRITE REGISTERS
  /////////////////////////////////


  //Write only register, clear on write (i.e. event)
  always @(posedge clk) begin
    if (!resetn_sync) begin
      reset_reg <= #1 `REG_RESET_DEFAULT;
    end else begin
      if (reg_wren) begin
        case (axi_awaddr)
          //Reset Register
          `REG_RESET_ADDR: begin
            for (
                byte_index = 0;
                byte_index <= (`REG_RESET_WIDTH / 8 - 1);
                byte_index = byte_index + 1
            )
            if (S_AXI_WSTRB[byte_index] == 1) begin
              reset_reg[byte_index*8+:8] <= S_AXI_WDATA[byte_index*8+:8];
            end
          end
          default: ;
        endcase
      end else begin
        reset_reg <= #1 `REG_RESET_DEFAULT;
      end
    end
  end

  //R/W register, not cleared
  always @(posedge clk) begin
    if (!resetn_sync) begin
      cpu2ip_flip_reg       <= #1 `REG_FLIP_DEFAULT;
      cpu2ip_debug_reg      <= #1 `REG_DEBUG_DEFAULT;
      cpu2ip_tgtipaddr_reg  <= #1 `REG_TGTIPADDR_DEFAULT;
      cpu2ip_tgtudpport_reg <= #1 `REG_TGTUDPPORT_DEFAULT;
    end else begin
      if (reg_wren)  //write event
        case (axi_awaddr)
          //Flip Register
          `REG_FLIP_ADDR: begin
            for (
                byte_index = 0; byte_index <= (`REG_FLIP_WIDTH / 8 - 1); byte_index = byte_index + 1
            )
            if (S_AXI_WSTRB[byte_index] == 1) begin  //dynamic register;
              cpu2ip_flip_reg[byte_index*8+:8] <= S_AXI_WDATA[byte_index*8+:8];
            end
          end
          //Debug Register
          `REG_DEBUG_ADDR: begin
            for (
                byte_index = 0;
                byte_index <= (`REG_DEBUG_WIDTH / 8 - 1);
                byte_index = byte_index + 1
            )
            if (S_AXI_WSTRB[byte_index] == 1) begin  // dynamic register;
              cpu2ip_debug_reg[byte_index*8+:8] <= S_AXI_WDATA[byte_index*8+:8];
            end
          end
          `REG_TGTIPADDR_ADDR: begin
            for (
                byte_index = 0;
                byte_index <= (`REG_TGTIPADDR_WIDTH / 8 - 1);
                byte_index = byte_index + 1
            )
            if (S_AXI_WSTRB[byte_index] == 1)  // dynamic register;
              cpu2ip_tgtipaddr_reg[byte_index*8+:8] <= S_AXI_WDATA[byte_index*8+:8];
          end
          `REG_TGTUDPPORT_ADDR: begin
            for (
                byte_index = 0;
                byte_index <= (`REG_TGTUDPPORT_WIDTH / 8 - 1);
                byte_index = byte_index + 1
            )
            if (S_AXI_WSTRB[byte_index] == 1)  // dynamic register;
              cpu2ip_tgtudpport_reg[byte_index*8+:8] <= S_AXI_WDATA[byte_index*8+:8];
          end
          default: ;
        endcase
    end
  end


  /////////////////////////////////
  ////    READ REGISTERS
  /////////////////////////////////


  // Implement memory mapped register select and read logic generation
  // Slave register read enable is asserted when valid address is available
  // and the slave is ready to accept the read address.

  // reg_rden control logic
  // temperary no extra logic here
  assign reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;

  always_comb begin
    case (axi_araddr)  // S_AXI_ARADDR ^ C_BASE_ADDRESS
      `REG_ID_ADDR:          reg_data_out[`REG_ID_BITS] = id_reg;
      `REG_VERSION_ADDR:     reg_data_out[`REG_VERSION_BITS] = version_reg;
      `REG_FLIP_ADDR:        reg_data_out[`REG_FLIP_BITS] = ip2cpu_flip_reg;
      `REG_DEBUG_ADDR:       reg_data_out[`REG_DEBUG_BITS] = ip2cpu_debug_reg;
      `REG_PKTIN_ADDR:       reg_data_out[`REG_PKTIN_BITS] = pktin_reg;
      `REG_PKTOUT_ADDR:      reg_data_out[`REG_PKTOUT_BITS] = pktout_reg;
      `REG_ICMPOUT_ADDR:     reg_data_out[`REG_ICMPOUT_BITS] = icmpout_reg;
      `REG_TGTIPADDR_ADDR:   reg_data_out[`REG_TGTIPADDR_BITS] = ip2cpu_tgtipaddr_reg;
      `REG_TGTIPOUT_ADDR:    reg_data_out[`REG_TGTIPOUT_BITS] = tgtipout_reg;
      `REG_TGTIPOUTLST_ADDR: reg_data_out[`REG_TGTIPOUTLST_BITS] = tgtipoutlst_reg;
      `REG_TGTUDPPORT_ADDR:  reg_data_out[`REG_TGTUDPPORT_BITS] = ip2cpu_tgtudpport_reg;
      `REG_TGTUDPCNT_ADDR:   reg_data_out[`REG_TGTUDPCNT_BITS] = tgtudpcnt_reg;
      default:               reg_data_out[31:0] = 32'hFEE1DEAD;  //Default return value
    endcase
  end  // end of assigning data to IP2Bus_Data bus

  // Read only registers, not cleared
  // Nothing to do here....

  // Read only registers, cleared on read (e.g. counters)
  always @(posedge clk)
    if (!resetn_sync) begin
      pktin_reg_clear      <= #1 1'b0;
      pktin_reg_clear_d    <= #1 1'b0;
      pktout_reg_clear     <= #1 1'b0;
      pktout_reg_clear_d   <= #1 1'b0;
      icmpout_reg_clear    <= #1 1'b0;
      icmpout_reg_clear_d  <= #1 1'b0;
      tgtipout_reg_clear   <= #1 1'b0;
      tgtipout_reg_clear_d <= #1 1'b0;
    end else begin
      pktin_reg_clear <= #1 pktin_reg_clear_d;
      pktin_reg_clear_d <= #1 (reg_rden && (axi_araddr == `REG_PKTIN_ADDR)) ? 1'b1 : 1'b0;
      pktout_reg_clear <= #1 pktout_reg_clear_d;
      pktout_reg_clear_d <= #1 (reg_rden && (axi_araddr == `REG_PKTOUT_ADDR)) ? 1'b1 : 1'b0;
      icmpout_reg_clear <= #1 icmpout_reg_clear_d;
      icmpout_reg_clear_d <= #1 (reg_rden && (axi_araddr == `REG_ICMPOUT_ADDR)) ? 1'b1 : 1'b0;
      tgtipout_reg_clear <= #1 tgtipout_reg_clear_d;
      tgtipout_reg_clear_d <= #1 (reg_rden && (axi_araddr == `REG_TGTIPOUT_ADDR)) ? 1'b1 : 1'b0;
    end


  // Output register or memory read data
  always @(posedge S_AXI_ACLK) begin
    if (S_AXI_ARESETN == 1'b0) begin
      axi_rdata <= 0;
    end else begin
      // When there is a valid read address (S_AXI_ARVALID) with
      // acceptance of read address by the slave (axi_arready),
      // output the read dada
      if (reg_rden) begin
        axi_rdata <= reg_data_out;  /*ip2bus_data*/  // register read data
      end
    end
  end
endmodule
